/***********************************************************
 * @author		Jon Hourany
 * @date		3/09/13
 * @class		EECE 444
 *
 * @file		ctrl_lines.v
 * @proj		Video Card
 ************************************************************/
module Top(RESET, H_SYNC, V_SYNC, RED, osc_clk);
	input  wire RESET;
	output wire H_SYNC;
	output wire V_SYNC;
	output wire RED;
	output wire osc_clk;
	//output reg  BLUE;	//output reg  GREEN;
	//output wire CLK_OUT;
	
	//event reset_trigger; 
     //event  reset_done_trigger; 
       
     //initial begin 
       //forever begin 
         //@ (reset_trigger); 
         //@ (negedge clk); 
         //reset = 0; 
         //@ (negedge clk); 
         //reset = 1; 
         //-> reset_done_trigger; 
       //end 
     //end
	 
	 //reg clk, reset;
	 //initial begin
		 //#1 reset 	= 0;
		 //#1 clk 	= 0;
		 //#2 reset 	= 1;
	 //end
	 
	 //always #1 clk = ~clk;
	//wire clk; 

	OSCC OSCC_1 (.OSC(osc_clk));
	CtrlLines CONTROLLINES(.NRST(reset), .CLK(osc_clk), .H_SYNC(H_SYNC), .V_SYNC(V_SYNC));
	
	assign RED = 1; 

	
endmodule 
